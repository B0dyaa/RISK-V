module Data_Mem(input clk,WE,input [31:0] WD,A,output reg [31:0] RD);
reg[7:0] Mem [31:0];
always @(posedge) begin
    
end
endmodule
